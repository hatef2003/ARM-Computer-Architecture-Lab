module IF (input clk , rst , branchTaken ,freeze ,input[31:0] branchAdrress ,output [31:0] PC,instruction )
    
endmodule;
