module memReg(input clk, rst, WB_EN ,MEM_R_EN ,input [31:0] AluRes ,input [3:0]dest);

endmodule