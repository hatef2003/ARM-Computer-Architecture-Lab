module IF_Reg(  input clk, rst, freeze, flush,
                input [31:0] pcIn, instructionIn,
                output reg [31:0] pc, Instruction);

endmodule